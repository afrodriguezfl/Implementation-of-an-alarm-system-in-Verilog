module Security_System()

endmodule 