module Security_System()

	always @(posedge clk)begin
	
	printf(Hola mundo);
	
	end
	
endmodule 