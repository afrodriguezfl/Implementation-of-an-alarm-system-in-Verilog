module Hola ()

endmodule
