`timescale 1ns / 1ps
module LCD_Top
(

		input CLOCK_50,       //50 MHz
		inout [7:0] LCD_DATA, //LCD Data bus 8 bits
		input [1:0] MESG,     //Message control signal
		output LCD_RW,        //LCD Read/Write Select, 0 = Write, 1 = Read
		output LCD_EN,        //LCD Enable
		output LCD_RS		    //LCD Command/Data Select, 0 = Command, 1 = Data

);

	reg [8:0] Mostrar_10  = "P";
	reg [8:0] Mostrar_11  = "R";
	reg [8:0] Mostrar_12  = "U";
	reg [8:0] Mostrar_13  = "E";
	reg [8:0] Mostrar_14  = "B";
	reg [8:0] Mostrar_15  = "A";
	reg [8:0] Mostrar_16  = " ";
	reg [8:0] Mostrar_17  = "L";
	reg [8:0] Mostrar_18  = "I";
	reg [8:0] Mostrar_19  = "N";
	reg [8:0] Mostrar_110 = "E";
	reg [8:0] Mostrar_111 = "A";
	reg [8:0] Mostrar_112 = " ";
	reg [8:0] Mostrar_113 = "1";
	reg [8:0] Mostrar_114 = " ";
	reg [8:0] Mostrar_115 = " ";
	reg [8:0] Mostrar_20  = "P";
	reg [8:0] Mostrar_21  = "R";
	reg [8:0] Mostrar_22  = "U";
	reg [8:0] Mostrar_23  = "E";
	reg [8:0] Mostrar_24  = "B";
	reg [8:0] Mostrar_25  = "A";
	reg [8:0] Mostrar_26  = " ";
	reg [8:0] Mostrar_27  = "L";
	reg [8:0] Mostrar_28  = "I";
	reg [8:0] Mostrar_29  = "N";
	reg [8:0] Mostrar_210 = "E";
	reg [8:0] Mostrar_211 = "A";
	reg [8:0] Mostrar_212 = " ";
	reg [8:0] Mostrar_213 = "2";
	reg [8:0] Mostrar_214 = " ";
	reg [8:0] Mostrar_215 = " ";               

	wire DLY_RST;

	Reset_Delay rst(.iCLK(CLOCK_50),.oRESET(DLY_RST));

	always @(CLOCK_50)begin

		case(MESG)

			0 : begin
				Mostrar_10  <= 9'h120;//Space
				Mostrar_11  <= 9'h153;//S
				Mostrar_12  <= 9'h154;//T
				Mostrar_13  <= 9'h141;//A
				Mostrar_14  <= 9'h154;//T
				Mostrar_15  <= 9'h155;//U
				Mostrar_16  <= 9'h153;//S
				Mostrar_17  <= 9'h13A;//:
				Mostrar_18  <= 9'h120;//Space
				Mostrar_19  <= 9'h16F;//o
				Mostrar_110 <= 9'h166;//f
				Mostrar_111 <= 9'h166;//f
				Mostrar_112 <= 9'h120;//Space
				Mostrar_113 <= 9'h120;//Space
				Mostrar_114 <= 9'h120;//Space
				Mostrar_115 <= 9'h120;//Space
				Mostrar_20  <= 9'h120;//Space
				Mostrar_21  <= 9'h157;//W
				Mostrar_22  <= 9'h13A;//:
				Mostrar_23  <= 9'h16E;//n
				Mostrar_24  <= 9'h16F;//o
				Mostrar_25  <= 9'h120;//Space
				Mostrar_26  <= 9'h153;//S
				Mostrar_27  <= 9'h13A;//:
				Mostrar_28  <= 9'h16E;//n
				Mostrar_29  <= 9'h16F;//o
				Mostrar_210 <= 9'h120; //Space
				Mostrar_211 <= 9'h14C;//L
				Mostrar_212 <= 9'h13A;//:
				Mostrar_213 <= 9'h16E;//n
				Mostrar_214 <= 9'h16F;//o
				Mostrar_215 <= 9'h120;//Space
			end

			1 : begin
				Mostrar_10  <= 9'h120;//Space
				Mostrar_11  <= 9'h153;//S
				Mostrar_12  <= 9'h154;//T
				Mostrar_13  <= 9'h141;//A
				Mostrar_14  <= 9'h154;//T
				Mostrar_15  <= 9'h155;//U
				Mostrar_16  <= 9'h153;//S
				Mostrar_17  <= 9'h13A;//:
				Mostrar_18  <= 9'h120;//Space
				Mostrar_19  <= 9'h16F;//o
				Mostrar_110 <= 9'h16e;//n
				Mostrar_111 <= 9'h120;//Space
				Mostrar_112 <= 9'h120;//Space
				Mostrar_113 <= 9'h120;//Space
				Mostrar_114 <= 9'h120;//Space
				Mostrar_115 <= 9'h120;//Space
				Mostrar_20  <= 9'h120;//Space
				Mostrar_21  <= 9'h157;//W
				Mostrar_22  <= 9'h13A;//:
				Mostrar_23  <= 9'h16E;//n
				Mostrar_24  <= 9'h16F;//o
				Mostrar_25  <= 9'h120;//Space
				Mostrar_26  <= 9'h153;//S
				Mostrar_27  <= 9'h13A;//:
				Mostrar_28  <= 9'h16E;//n
				Mostrar_29  <= 9'h16F;//o
				Mostrar_210 <= 9'h120; //Space
				Mostrar_211 <= 9'h14C;//L
				Mostrar_212 <= 9'h13A;//:
				Mostrar_213 <= 9'h16E;//n
				Mostrar_214 <= 9'h16F;//o
				Mostrar_215 <= 9'h120;//Space
				end
				
			2 : begin
				Mostrar_10  <= 9'h120;//Space
				Mostrar_11  <= 9'h153;//S
				Mostrar_12  <= 9'h154;//T
				Mostrar_13  <= 9'h141;//A
				Mostrar_14  <= 9'h154;//T
				Mostrar_15  <= 9'h155;//U
				Mostrar_16  <= 9'h153;//S
				Mostrar_17  <= 9'h13A;//:
				Mostrar_18  <= 9'h120;//Space
				Mostrar_19  <= 9'h161;//a
				Mostrar_110 <= 9'h16C;//l
				Mostrar_111 <= 9'h161;//a
				Mostrar_112 <= 9'h172;//r
				Mostrar_113 <= 9'h16D;//m
				Mostrar_114 <= 9'h120;//Space
				Mostrar_115 <= 9'h120;//Space
				Mostrar_20  <= 9'h120;//Space
				Mostrar_21  <= 9'h157;//W
				Mostrar_22  <= 9'h13A;//:
				Mostrar_23  <= 9'h173;//s
				Mostrar_24  <= 9'h169;//i
				Mostrar_25  <= 9'h120;//Space
				Mostrar_26  <= 9'h153;//S
				Mostrar_27  <= 9'h13A;//:
				Mostrar_28  <= 9'h173;//s
				Mostrar_29  <= 9'h169;//i
				Mostrar_210 <= 9'h120; //Space
				Mostrar_211 <= 9'h14C;//L
				Mostrar_212 <= 9'h13A;//:
				Mostrar_213 <= 9'h16E;//n
				Mostrar_214 <= 9'h16F;//o
				Mostrar_215 <= 9'h120;//Space
			end
			
			3 : begin
				Mostrar_10  <= 9'h120;//Space
				Mostrar_11  <= 9'h153;//S
				Mostrar_12  <= 9'h154;//T
				Mostrar_13  <= 9'h141;//A
				Mostrar_14  <= 9'h154;//T
				Mostrar_15  <= 9'h155;//U
				Mostrar_16  <= 9'h153;//S
				Mostrar_17  <= 9'h13A;//:
				Mostrar_18  <= 9'h120;//Space
				Mostrar_19  <= 9'h164;//d
				Mostrar_110 <= 9'h161;//a
				Mostrar_111 <= 9'h16E;//n
				Mostrar_112 <= 9'h167;//g
				Mostrar_113 <= 9'h165;//e
				Mostrar_114 <= 9'h172;//r
				Mostrar_115 <= 9'h120;//Space
				Mostrar_20  <= 9'h120;//Space
				Mostrar_21  <= 9'h157;//W
				Mostrar_22  <= 9'h13A;//:
				Mostrar_23  <= 9'h173;//s
				Mostrar_24  <= 9'h169;//i
				Mostrar_25  <= 9'h120;//Space
				Mostrar_26  <= 9'h153;//S
				Mostrar_27  <= 9'h13A;//:
				Mostrar_28  <= 9'h173;//s
				Mostrar_29  <= 9'h169;//i
				Mostrar_210 <= 9'h120; //Space
				Mostrar_211 <= 9'h14C;//L
				Mostrar_212 <= 9'h13A;//:
				Mostrar_213 <= 9'h173;//s
				Mostrar_214 <= 9'h169;//i
				Mostrar_215 <= 9'h120;//Space
			end

		endcase

	end

	LCD_Write wrt(
	
	/////////////HOST SIDE//////////////////
		.iCLK(CLOCK_50),
		.iRST_N(DLY_RST),
	////////////////////////////////////////
	
	//////////////LCD SIDE//////////////////
		.LCD_DATA(LCD_DATA),
		.LCD_RW(LCD_RW),
		.LCD_EN(LCD_EN),
		.LCD_RS(LCD_RS),   
		.Mostrar_10(Mostrar_10),
		.Mostrar_11(Mostrar_11),
		.Mostrar_12(Mostrar_12),
		.Mostrar_13(Mostrar_13),
		.Mostrar_14(Mostrar_14),
		.Mostrar_15(Mostrar_15),
		.Mostrar_16(Mostrar_16),
		.Mostrar_17(Mostrar_17),
		.Mostrar_18(Mostrar_18),
		.Mostrar_19(Mostrar_19),
		.Mostrar_110(Mostrar_110),
		.Mostrar_111(Mostrar_111),
		.Mostrar_112(Mostrar_112),
		.Mostrar_113(Mostrar_113),
		.Mostrar_114(Mostrar_114),
		.Mostrar_115(Mostrar_115),
		.Mostrar_20(Mostrar_20),
		.Mostrar_21(Mostrar_21),
		.Mostrar_22(Mostrar_22),
		.Mostrar_23(Mostrar_23),
		.Mostrar_24(Mostrar_24),
		.Mostrar_25(Mostrar_25),
		.Mostrar_26(Mostrar_26),
		.Mostrar_27(Mostrar_27),
		.Mostrar_28(Mostrar_28),
		.Mostrar_29(Mostrar_29),
		.Mostrar_210(Mostrar_210),
		.Mostrar_211(Mostrar_211),
		.Mostrar_212(Mostrar_212),
		.Mostrar_213(Mostrar_213),
		.Mostrar_214(Mostrar_214),
		.Mostrar_215(Mostrar_215)
	////////////////////////////////////////
	
);

endmodule
